-- A DUT entity is used to wrap your design.
--  This example shows how you can do this for the
--  Full-adder.

library ieee;
use ieee.std_logic_1164.all;

entity DUT is
   port(input_vector: in std_logic_vector(127 downto 0);
       	output_vector: out std_logic_vector(1407 downto 0));
end entity;

architecture DutWrap of DUT is
	-- Instantiate your own top Module component in place of ALU_1
	Component keyexp is
	port (key: in std_logic_vector(127 downto 0); outp:out std_logic_vector (1407 downto 0));
	end component keyexp;
begin

   -- input/output vector element ordering is critical,
   -- and must match the ordering in the trace file!
   add_instance: keyexp port map (key => input_vector(127 downto 0), outp => output_vector(1407 downto 0));

end DutWrap;